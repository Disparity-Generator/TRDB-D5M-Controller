-- megafunction wizard: %LPM_DIVIDE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_DIVIDE 

-- ============================================================
-- File Name: Teiler_12_Bit.vhd
-- Megafunction Name(s):
-- 			LPM_DIVIDE
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2020  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.all;

ENTITY Teiler_12_Bit IS
	PORT
	(
		denom		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		numer		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		quotient		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
		remain		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0)
	);
END Teiler_12_Bit;


ARCHITECTURE SYN OF teiler_12_bit IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (11 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (11 DOWNTO 0);



	COMPONENT lpm_divide
	GENERIC (
		lpm_drepresentation		: STRING;
		lpm_hint		: STRING;
		lpm_nrepresentation		: STRING;
		lpm_type		: STRING;
		lpm_widthd		: NATURAL;
		lpm_widthn		: NATURAL
	);
	PORT (
			denom	: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			numer	: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			quotient	: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			remain	: OUT STD_LOGIC_VECTOR (11 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	quotient    <= sub_wire0(11 DOWNTO 0);
	remain    <= sub_wire1(11 DOWNTO 0);

	LPM_DIVIDE_component : LPM_DIVIDE
	GENERIC MAP (
		lpm_drepresentation => "UNSIGNED",
		lpm_hint => "LPM_REMAINDERPOSITIVE=TRUE",
		lpm_nrepresentation => "UNSIGNED",
		lpm_type => "LPM_DIVIDE",
		lpm_widthd => 12,
		lpm_widthn => 12
	)
	PORT MAP (
		denom => denom,
		numer => numer,
		quotient => sub_wire0,
		remain => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
-- Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
-- Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "0"
-- Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE"
-- Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
-- Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "12"
-- Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "12"
-- Retrieval info: USED_PORT: denom 0 0 12 0 INPUT NODEFVAL "denom[11..0]"
-- Retrieval info: USED_PORT: numer 0 0 12 0 INPUT NODEFVAL "numer[11..0]"
-- Retrieval info: USED_PORT: quotient 0 0 12 0 OUTPUT NODEFVAL "quotient[11..0]"
-- Retrieval info: USED_PORT: remain 0 0 12 0 OUTPUT NODEFVAL "remain[11..0]"
-- Retrieval info: CONNECT: @denom 0 0 12 0 denom 0 0 12 0
-- Retrieval info: CONNECT: @numer 0 0 12 0 numer 0 0 12 0
-- Retrieval info: CONNECT: quotient 0 0 12 0 @quotient 0 0 12 0
-- Retrieval info: CONNECT: remain 0 0 12 0 @remain 0 0 12 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Teiler_12_Bit.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Teiler_12_Bit.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Teiler_12_Bit.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Teiler_12_Bit.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Teiler_12_Bit_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
